/// # guid

/// ## guid

/// ### guid
nominal guid_python =
    `(
        global "import uuid"
        $'' : $'uuid.UUID'
    )
type guid_switch =
    {
        Fsharp : $'System.Guid'
        Python : guid_python
    }
nominal guid = $'backend_switch `(guid_switch)'

/// ### new_guid
inl new_guid (x : string) : guid =
    run_target_args (fun () => x) function
        | Rust (Contract) => fun _ => null ()
        | _ => fun x => x |> convert

/// ### new_raw_guid
inl new_raw_guid () : guid =
    backend_switch {
        Fsharp = fun () => $'System.Guid.NewGuid' () : guid
        Python = fun () => $'uuid.uuid4()' : guid
    }

/// ### hash_guid
type hash_guid = guid

let hash_guid (hash : string) : hash_guid =
    inl hash = hash |> sm'.pad_left 32i32 '0'
    run_target_args (fun () => hash) function
        | Rust (Contract) => fun _ => null ()
        | _ => fun hash =>
            inl a = hash |> sm'.range (am'.Start 0i32) (am'.End fun _ => 8)
            inl b = hash |> sm'.range (am'.Start 8i32) (am'.End fun _ => 12)
            inl c = hash |> sm'.range (am'.Start 12i32) (am'.End fun _ => 16)
            inl d = hash |> sm'.range (am'.Start 16i32) (am'.End fun _ => 20)
            inl e = hash |> sm'.range (am'.Start 20i32) (am'.End fun _ => 32)
            $'$"{!a}-{!b}-{!c}-{!d}-{!e}"' |> new_guid

/// ## main
inl main () =
    $'let new_guid x = !new_guid x' : ()
    $'let hash_guid x = !hash_guid x' : ()
    $'let new_raw_guid x = !new_raw_guid x' : ()
