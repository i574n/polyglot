open rust_operators

inl main (args : array_base string) =
    leptos.log $'"main / args: " + string !args + ""'

    !\($'"let _ = console_log::init_with_level(log::Level::Debug)"')
    !\($'"console_error_panic_hook::set_once()"')

    inl body : optionm'.option' rust.html_element = !\($'"leptos::document().body()"')
    inl body = body |> optionm'.unbox
    inl body_log = body |> sm'.format_debug

    leptos.log $'"main / mount_to_body / body: " + string !body_log + ""'

    let mount () =
        fun () =>
            src.components.app.render ()
            |> leptos.to_view_trait
        |> leptos.mount_to_body

    match body with
    | Some body =>
        body |> leptos.set_inner_html ""

        mount ()
    | _ =>
        inl fn : rust.box (rust.dyn' rust.fn_unit) = rust.box_fn mount
        inl fn_closure = fn |> rust.closure_wrap
        inl fn = fn_closure |> rust.closure_as_ref |> rust.unchecked_ref

        !\($'"leptos::document().add_event_listener_with_callback(\\\"DOMContentLoaded\\\", !fn).unwrap()"')

        fn_closure |> rust.closure_forget

    0i32

inl main () =
    print_static "<dice_ui>"
    rust.types ()
    leptos.types ()
    src.model.near.backend.types ()

    $"let main args = !main args" : ()
    print_static "</dice_ui>"
