/// # parsing
open rust_operators
open sm'_operators

/// ## types
inl types () =
    ()

inl types () =
    types ()

/// ## fparsec

/// ## range
type range =
    {
        from : int
        to : int
    }

/// ## position
type position =
    {
        line : int
        col : int
    }

/// ## parser_state
type parser_state =
    {
        line_text : sm'.string_builder
        position : position
    }

/// ## parser
type parser t = string * parser_state -> result (t * string * parser_state) string

/// ## parse
inl parse forall t. (p : parser t) (input : string) : result (t * string * parser_state) string =
    p (input, { line_text = "" |> sm'.string_builder; position = { line = 1; col = 1 } })

/// ## inc
inl inc c (s : parser_state) =
    match c with
    | '\n' => { line = s.position.line + 1; col = 1 }
    | _ => { s.position with col = s.position.col + 1 }.position

/// ## update
inl update result (s : parser_state) =
    (s, result |> sm'.to_char_array |> am'.to_list' |> listm'.unbox)
    ||> listm.fold fun s c => { s with
        position = s |> inc c
        line_text =
            match c with
            | '\n' => s.line_text |> sm'.builder_clear
            | c => s.line_text |> sm'.builder_append (sm'.obj_to_string c)
    }

/// ## any_char
inl any_char () : parser char = function
    | "", s => Error $'$"parsing.any_char / unexpected end of input / s: %A{!s}"'
    | x, s =>
        inl first_char = x |> sm'.index 0i32
        inl rest = x |> sm'.range (am'.Start 1i32) (am'.End id)
        in Ok (first_char, rest, s |> update (sm'.obj_to_string first_char))

/// ## p_char
inl p_char (c : char) : parser char = function
    | "", s => Error $'$"parsing.p_char / unexpected end of input / s: %A{!s}"'
    | input, s =>
        inl first_char = input |> sm'.index 0i32
        if first_char = c
        then Ok (
            first_char,
            input |> sm'.range (am'.Start 1i32) (am'.End id),
            s |> update (sm'.obj_to_string first_char)
        )
        else
            inl { line_text position = { line col } } = s
            inl message : string =
                inl rest =
                    input
                    |> sm'.range
                        (am'.Start 0i32)
                        (am'.End fun l =>
                            match (input |> sm'.index_of "\n") - 1 with
                            | -2 => l
                            | l => l
                        )
                $'$"parsing.p_char / expected: \'{!c}\' / line: {!line} / col: {!col}\n{!line_text}{!rest}"'
            inl pointer_line = (sm'.replicate (col - 1) " ") +. "^"
            $'$"{!message}\n{!pointer_line}\n"' |> Error

/// ## any_string
inl any_string length : parser string = fun input, s =>
    if sm'.length input < length
    then Error $'$"parsing.any_string / unexpected end of input / s: %A{!s}"'
    else
        inl result = input |> sm'.range (am'.Start 0i32) (am'.End fun _ => length - 1)
        inl rest = input |> sm'.range (am'.Start length) (am'.End id)
        Ok (result, rest, s |> update result)

/// ## skip_any_string
inl skip_any_string length : parser () = fun input, s =>
    if sm'.length input < length
    then Error $'$"parsing.skip_any_string / unexpected end of input / s: %A{!s}"'
    else Ok (
        (),
        input |> sm'.range (am'.Start length) (am'.End id),
        s |> update (input |> sm'.range (am'.Start 0i32) (am'.End fun _ => length - 1))
    )

/// ## (>>.)
inl (>>.) forall t u. (a : parser t) (b : parser u) : parser u = fun input, s =>
    match a (input, s) with
    | Ok (_, rest, s) => b (rest, s)
    | Error e => Error e

/// ## none_of
inl none_of (chars : list char) : parser char = function
    | "", s =>
        inl chars = chars |> listm'.box |> listm'.to_array'
        Error $'$"parsing.none_of / unexpected end of input / chars: %A{!chars} / s: %A{!s}"'
    | x, s =>
        inl first_char = x |> sm'.index 0i32
        inl rest = x |> sm'.range (am'.Start 1i32) (am'.End id)
        if chars |> listm'.exists' ((=) first_char) |> not
        then Ok (first_char, rest, s |> update (sm'.obj_to_string first_char))
        else
            inl chars = chars |> listm'.box |> listm'.to_array'
            Error $'$"parsing.none_of / unexpected char: \'{!first_char}\' / chars: %A{!chars} / s: %A{!s}"'

/// ## (<|>)
inl (<|>) forall t. (a : parser t) (b : parser t) : parser t = fun input, s =>
    match a (input, s) with
    | Ok _ as result => result
    | Error _ => b (input, s)

/// ## (|>>)
inl (|>>) p f : parser _ = fun input =>
    match p input with
    | Ok (result, rest) => Ok (f result, rest)
    | Error e => Error e

/// ## many1_chars
inl many1_chars p : parser string = fun input =>
    match p input with
    | Error e => Error e
    | Ok (first_result, rest) =>
        let rec loop acc input =
            match p input with
            | Ok (result, rest) => loop (acc +. sm'.obj_to_string result) rest
            | Error _ => Ok (acc, input)
        loop (sm'.obj_to_string first_result) rest

/// ## many1
inl many1 p : parser (list _) = fun input =>
    match p input with
    | Error e => Error e
    | Ok (first_result, rest) =>
        let rec loop acc input =
            match p input with
            | Ok (result, rest) => loop (result :: acc) rest
            | Error _ => Ok (listm.rev acc, input)
        loop [ first_result ] rest

/// ## many1_strings
inl many1_strings p : parser string = fun input =>
    match many1 p input with
    | Ok (results, rest) =>
        Ok (results |> listm.map sm'.obj_to_string |> listm'.box |> seq.of_list' |> sm'.concat "", rest)
    | Error e => Error e

/// ## choice
inl choice parsers : parser _ = fun input =>
    let rec loop = function
        | [] => Error "choice / no parsers succeeded"
        | p :: ps =>
            match p input with
            | Ok _ as result => result
            | Error _ => loop ps
    loop parsers

/// ## many
inl many p : parser (list _) = fun input =>
    let rec loop acc input =
        match p input with
        | Ok (result, rest) => loop (result :: acc) rest
        | Error _ => Ok (listm.rev acc, input)
    loop [] input

/// ## between
inl between p_open p_close p_content : parser _ = fun input =>
    match p_open input with
    | Ok (_, rest1) =>
        match p_content rest1 with
        | Ok (result, rest2) =>
            match p_close rest2 with
            | Ok (_, rest3) => Ok (result, rest3)
            | Error e => Error $'$"between / expected closing delimiter / e: %A{!e} / input: %A{!input} / rest1: %A{!rest1} / rest2: %A{!rest2}"'
        | Error _ => Error "between / expected content"
    | Error e => Error e

/// ## sep_by
inl sep_by p sep : parser (list _) = fun input, s =>
    let rec loop acc input s =
        match p (input, s) with
        | Error _ => Ok (acc |> listm.rev, input, s)
        | Ok (result, rest, s) =>
            match sep (rest, s) with
            | Error _ => Ok ((result :: acc) |> listm.rev, rest, s)
            | Ok (_, rest, s) => loop (result :: acc) rest s
    loop [] input s

/// ## span
inl span pred str =
    let rec loop i =
        if i >= sm'.length str
        then i
        elif pred (str |> sm'.index i)
        then loop (i + 1)
        else i
    loop 0

/// ## spaces1
inl spaces1 () : parser () = fun input, s =>
    match input |> span fun c => c = ' ' with
    | 0i32 => Error "spaces1 / expected at least one space"
    | n => Ok ((), input |> sm'.range (am'.Start n) (am'.End id), s)

/// ## p_digit
inl p_digit () : parser char = fun input, s =>
    match input |> sm'.index 0i32 with
    | ('0' | '1' | '2' | '3' | '4' | '5' | '6' | '7' | '8' | '9') as c =>
        Ok (c, input |> sm'.range (am'.Start 1i32) (am'.End id), s)
    | c => Error $'$"p_digit / unexpected char: {!c}"'
