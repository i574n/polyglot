/// # guid

/// ## guid

/// ### guid
nominal guid_python =
    `(
        global "import uuid"
        $'' : $'uuid.UUID'
    )
type guid_switch =
    {
        Fsharp : $'System.Guid'
        Python : guid_python
    }
nominal guid = $'backend_switch `(guid_switch)'

/// ### new_guid
inl new_guid (x : string) : guid =
    x |> convert

/// ### new_raw_guid
inl new_raw_guid () : guid =
    backend_switch {
        Fsharp = fun () => $'System.Guid.NewGuid' () : guid
        Python = fun () => $'uuid.uuid4()' : guid
    }

/// ### hash_guid
type hash_guid = guid

let hash_guid (~hash : string) : hash_guid =
    run_target function
        | Rust (Contract) => fun () => null ()
        | _ => fun () =>
            inl hash = hash |> sm'.pad_left 32i32 '0'
            inl a = hash |> sm'.range (am'.Start 0i32) (am'.End fun _ => 8)
            inl b = hash |> sm'.range (am'.Start 8i32) (am'.End fun _ => 12)
            inl c = hash |> sm'.range (am'.Start 12i32) (am'.End fun _ => 16)
            inl d = hash |> sm'.range (am'.Start 16i32) (am'.End fun _ => 20)
            inl e = hash |> sm'.range (am'.Start 20i32) (am'.End fun _ => 32)
            $'$"{!a}-{!b}-{!c}-{!d}-{!e}"' : string
            |> fun x => x : string
            |> convert

/// ## main
inl main () =
    $'let new_guid x = !new_guid x' : ()
    $'let hash_guid x = !hash_guid x' : ()
    $'let new_raw_guid x = !new_raw_guid x' : ()
